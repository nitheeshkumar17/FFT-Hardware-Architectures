`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:06:34 07/18/2019 
// Design Name: 
// Module Name:    buf_25 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module buf_25(
    input [31:0] a_re,
    input [31:0] a_img,
    input [31:0] b_re,
    input [31:0] b_img,
    input clk,
    output reg [31:0] a1_re,
    output reg [31:0] a1_img,
    output reg [31:0] b1_re,
    output reg [31:0] b1_img
    );

reg [31:0] n0 [0:26];
reg [31:0] n1 [0:26];
reg [31:0] n2 [0:26];
reg [31:0] n3 [0:26];
always @(posedge clk) begin
n0[0]<=a_re;
n0[1]<=n0[0];
n0[2]<=n0[1];
n0[3]<=n0[2];
n0[4]<=n0[3];
n0[5]<=n0[4];
n0[6]<=n0[5];
n0[7]<=n0[6];
n0[8]<=n0[7];
n0[9]<=n0[8];
n0[10]<=n0[9];
n0[11]<=n0[10];
n0[12]<=n0[11];
n0[13]<=n0[12];
n0[14]<=n0[13];
n0[15]<=n0[14];
n0[16]<=n0[15];
n0[17]<=n0[16];
n0[18]<=n0[17];
n0[19]<=n0[18];
n0[20]<=n0[19];
n0[21]<=n0[20];
n0[22]<=n0[21];
n0[23]<=n0[22];
n0[24]<=n0[23];
n0[25]<=n0[24];
n0[26]<=n0[25];
a1_re<=n0[26];


n1[0]<=a_img;
n1[1]<=n1[0];
n1[2]<=n1[1];
n1[3]<=n1[2];
n1[4]<=n1[3];
n1[5]<=n1[4];
n1[6]<=n1[5];
n1[7]<=n1[6];
n1[8]<=n1[7];
n1[9]<=n1[8];
n1[10]<=n1[9];
n1[11]<=n1[10];
n1[12]<=n1[11];
n1[13]<=n1[12];
n1[14]<=n1[13];
n1[15]<=n1[14];
n1[16]<=n1[15];
n1[17]<=n1[16];
n1[18]<=n1[17];
n1[19]<=n1[18];
n1[20]<=n1[19];
n1[21]<=n1[20];
n1[22]<=n1[21];
n1[23]<=n1[22];
n1[24]<=n1[23];
n1[25]<=n1[24];
n1[26]<=n1[25];
a1_img<=n1[26];

n2[0]<=b_re;
n2[1]<=n2[0];
n2[2]<=n2[1];
n2[3]<=n2[2];
n2[4]<=n2[3];
n2[5]<=n2[4];
n2[6]<=n2[5];
n2[7]<=n2[6];
n2[8]<=n2[7];
n2[9]<=n2[8];
n2[10]<=n2[9];
n2[11]<=n2[10];
n2[12]<=n2[11];
n2[13]<=n2[12];
n2[14]<=n2[13];
n2[15]<=n2[14];
n2[16]<=n2[15];
n2[17]<=n2[16];
n2[18]<=n2[17];
n2[19]<=n2[18];
n2[20]<=n2[19];
n2[21]<=n2[20];
n2[22]<=n2[21];
n2[23]<=n2[22];
n2[24]<=n2[23];
n2[25]<=n2[24];
n2[26]<=n2[25];
b1_re<=n2[26];

n3[0]<=b_img;
n3[1]<=n3[0];
n3[2]<=n3[1];
n3[3]<=n3[2];
n3[4]<=n3[3];
n3[5]<=n3[4];
n3[6]<=n3[5];
n3[7]<=n3[6];
n3[8]<=n3[7];
n3[9]<=n3[8];
n3[10]<=n3[9];
n3[11]<=n3[10];
n3[12]<=n3[11];
n3[13]<=n3[12];
n3[14]<=n3[13];
n3[15]<=n3[14];
n3[16]<=n3[15];
n3[17]<=n3[16];
n3[18]<=n3[17];
n3[19]<=n3[18];
n3[20]<=n3[19];
n3[21]<=n3[20];
n3[22]<=n3[21];
n3[23]<=n3[22];
n3[24]<=n3[23];
n3[25]<=n3[24];
n3[26]<=n3[25];
b1_img<=n3[26];
end

endmodule
