`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:39:49 07/26/2019 
// Design Name: 
// Module Name:    buf_30 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module buf_30(
    input [31:0] a_re,
    input [31:0] a_img,
    input clk,
    output reg [31:0] a1_re,
    output reg [31:0] a1_img
    );

reg [31:0] n0 [0:28];
reg [31:0] n1 [0:28];
always @(posedge clk) begin
n0[0]<=a_re;
n0[1]<=n0[0];
n0[2]<=n0[1];
n0[3]<=n0[2];
n0[4]<=n0[3];
n0[5]<=n0[4];
n0[6]<=n0[5];
n0[7]<=n0[6];
n0[8]<=n0[7];
n0[9]<=n0[8];
n0[10]<=n0[9];
n0[11]<=n0[10];
n0[12]<=n0[11];
n0[13]<=n0[12];
n0[14]<=n0[13];
n0[15]<=n0[14];
n0[16]<=n0[15];
n0[17]<=n0[16];
n0[18]<=n0[17];
n0[19]<=n0[18];
n0[20]<=n0[19];
n0[21]<=n0[20];
n0[22]<=n0[21];
n0[23]<=n0[22];
n0[24]<=n0[23];
n0[25]<=n0[24];
n0[26]<=n0[25];
n0[27]<=n0[26];
n0[28]<=n0[27];
a1_re<=n0[28];

n1[0]<=a_img;
n1[1]<=n1[0];
n1[2]<=n1[1];
n1[3]<=n1[2];
n1[4]<=n1[3];
n1[5]<=n1[4];
n1[6]<=n1[5];
n1[7]<=n1[6];
n1[8]<=n1[7];
n1[9]<=n1[8];
n1[10]<=n1[9];
n1[11]<=n1[10];
n1[12]<=n1[11];
n1[13]<=n1[12];
n1[14]<=n1[13];
n1[15]<=n1[14];
n1[16]<=n1[15];
n1[17]<=n1[16];
n1[18]<=n1[17];
n1[19]<=n1[18];
n1[20]<=n1[19];
n1[21]<=n1[20];
n1[22]<=n1[21];
n1[23]<=n1[22];
n1[24]<=n1[23];
n1[25]<=n1[24];
n1[26]<=n1[25];
n1[27]<=n1[26];
n1[28]<=n1[27];
a1_img<=n1[28];
end

endmodule
